
`define BITS 64
`define PINS 16
`define STACK_DEPTH 16
`define STACK_PTR_WIDTH 4 
