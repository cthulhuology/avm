
`define BITS 16
`define PINS 16
`define DEPTH 16
`define PTR 4 
